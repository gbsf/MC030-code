include/common_cells/assertions.svh