include/common_cells/registers.svh